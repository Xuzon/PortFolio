----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    21:39:50 11/05/2015 
-- Design Name: 
-- Module Name:    consulta_luz - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity consulta_luz is
    Port ( dir_lut : in  STD_LOGIC_VECTOR (7 downto 0);
           luz_id : out  STD_LOGIC_VECTOR (7 downto 0));
end consulta_luz;

architecture Behavioral of consulta_luz is

begin

luz_id <= "00001000" WHEN dir_lut ="00000000" ELSE
"00010010" WHEN dir_lut ="00000001" ELSE
"00100100" WHEN dir_lut ="00000010" ELSE
"00101110" WHEN dir_lut ="00000011" ELSE
"01010101" WHEN dir_lut ="00000100" ELSE
"10000000" WHEN dir_lut ="00000101" ELSE
"10100000" WHEN dir_lut ="00000110" ELSE
"10100100" WHEN dir_lut ="00000111" ELSE
"10100111" WHEN dir_lut ="00001000" ELSE
"10101010" WHEN dir_lut ="00001001" ELSE
"10101101" WHEN dir_lut ="00001010" ELSE
"10101111" WHEN dir_lut ="00001011" ELSE
"10110001" WHEN dir_lut ="00001100" ELSE
"10110011" WHEN dir_lut ="00001101" ELSE
"10110101" WHEN dir_lut ="00001110" ELSE
"10110111" WHEN dir_lut ="00001111" ELSE
"10111001" WHEN dir_lut ="00010000" ELSE
"10111010" WHEN dir_lut ="00010001" ELSE
"10111100" WHEN dir_lut ="00010010" ELSE
"10111101" WHEN dir_lut ="00010011" ELSE
"10111110" WHEN dir_lut ="00010100" ELSE
"10111111" WHEN dir_lut ="00010101" ELSE
"11000001" WHEN dir_lut ="00010110" ELSE
"11000010" WHEN dir_lut ="00010111" ELSE
"11000011" WHEN dir_lut ="00011000" ELSE
"11000100" WHEN dir_lut ="00011001" ELSE
"11000101" WHEN dir_lut ="00011010" ELSE
"11000110" WHEN dir_lut ="00011011" ELSE
"11000111" WHEN dir_lut ="00011100" ELSE
"11001000" WHEN dir_lut ="00011101" ELSE
"11001000" WHEN dir_lut ="00011110" ELSE
"11001001" WHEN dir_lut ="00011111" ELSE
"11001010" WHEN dir_lut ="00100000" ELSE
"11001011" WHEN dir_lut ="00100001" ELSE
"11001100" WHEN dir_lut ="00100010" ELSE
"11001100" WHEN dir_lut ="00100011" ELSE
"11001101" WHEN dir_lut ="00100100" ELSE
"11001110" WHEN dir_lut ="00100101" ELSE
"11001110" WHEN dir_lut ="00100110" ELSE
"11001111" WHEN dir_lut ="00100111" ELSE
"11010000" WHEN dir_lut ="00101000" ELSE
"11010000" WHEN dir_lut ="00101001" ELSE
"11010001" WHEN dir_lut ="00101010" ELSE
"11010010" WHEN dir_lut ="00101011" ELSE
"11010010" WHEN dir_lut ="00101100" ELSE
"11010011" WHEN dir_lut ="00101101" ELSE
"11010011" WHEN dir_lut ="00101110" ELSE
"11010100" WHEN dir_lut ="00101111" ELSE
"11010100" WHEN dir_lut ="00110000" ELSE
"11010101" WHEN dir_lut ="00110001" ELSE
"11010101" WHEN dir_lut ="00110010" ELSE
"11010110" WHEN dir_lut ="00110011" ELSE
"11010110" WHEN dir_lut ="00110100" ELSE
"11010111" WHEN dir_lut ="00110101" ELSE
"11010111" WHEN dir_lut ="00110110" ELSE
"11011000" WHEN dir_lut ="00110111" ELSE
"11011000" WHEN dir_lut ="00111000" ELSE
"11011001" WHEN dir_lut ="00111001" ELSE
"11011001" WHEN dir_lut ="00111010" ELSE
"11011010" WHEN dir_lut ="00111011" ELSE
"11011010" WHEN dir_lut ="00111100" ELSE
"11011010" WHEN dir_lut ="00111101" ELSE
"11011011" WHEN dir_lut ="00111110" ELSE
"11011011" WHEN dir_lut ="00111111" ELSE
"11011100" WHEN dir_lut ="01000000" ELSE
"11011100" WHEN dir_lut ="01000001" ELSE
"11011100" WHEN dir_lut ="01000010" ELSE
"11011101" WHEN dir_lut ="01000011" ELSE
"11011101" WHEN dir_lut ="01000100" ELSE
"11011110" WHEN dir_lut ="01000101" ELSE
"11011110" WHEN dir_lut ="01000110" ELSE
"11011110" WHEN dir_lut ="01000111" ELSE
"11011111" WHEN dir_lut ="01001000" ELSE
"11011111" WHEN dir_lut ="01001001" ELSE
"11011111" WHEN dir_lut ="01001010" ELSE
"11100000" WHEN dir_lut ="01001011" ELSE
"11100000" WHEN dir_lut ="01001100" ELSE
"11100000" WHEN dir_lut ="01001101" ELSE
"11100001" WHEN dir_lut ="01001110" ELSE
"11100001" WHEN dir_lut ="01001111" ELSE
"11100001" WHEN dir_lut ="01010000" ELSE
"11100010" WHEN dir_lut ="01010001" ELSE
"11100010" WHEN dir_lut ="01010010" ELSE
"11100010" WHEN dir_lut ="01010011" ELSE
"11100011" WHEN dir_lut ="01010100" ELSE
"11100011" WHEN dir_lut ="01010101" ELSE
"11100011" WHEN dir_lut ="01010110" ELSE
"11100011" WHEN dir_lut ="01010111" ELSE
"11100100" WHEN dir_lut ="01011000" ELSE
"11100100" WHEN dir_lut ="01011001" ELSE
"11100100" WHEN dir_lut ="01011010" ELSE
"11100101" WHEN dir_lut ="01011011" ELSE
"11100101" WHEN dir_lut ="01011100" ELSE
"11100101" WHEN dir_lut ="01011101" ELSE
"11100101" WHEN dir_lut ="01011110" ELSE
"11100110" WHEN dir_lut ="01011111" ELSE
"11100110" WHEN dir_lut ="01100000" ELSE
"11100110" WHEN dir_lut ="01100001" ELSE
"11100110" WHEN dir_lut ="01100010" ELSE
"11100111" WHEN dir_lut ="01100011" ELSE
"11100111" WHEN dir_lut ="01100100" ELSE
"11100111" WHEN dir_lut ="01100101" ELSE
"11100111" WHEN dir_lut ="01100110" ELSE
"11101000" WHEN dir_lut ="01100111" ELSE
"11101000" WHEN dir_lut ="01101000" ELSE
"11101000" WHEN dir_lut ="01101001" ELSE
"11101000" WHEN dir_lut ="01101010" ELSE
"11101001" WHEN dir_lut ="01101011" ELSE
"11101001" WHEN dir_lut ="01101100" ELSE
"11101001" WHEN dir_lut ="01101101" ELSE
"11101001" WHEN dir_lut ="01101110" ELSE
"11101010" WHEN dir_lut ="01101111" ELSE
"11101010" WHEN dir_lut ="01110000" ELSE
"11101010" WHEN dir_lut ="01110001" ELSE
"11101010" WHEN dir_lut ="01110010" ELSE
"11101010" WHEN dir_lut ="01110011" ELSE
"11101011" WHEN dir_lut ="01110100" ELSE
"11101011" WHEN dir_lut ="01110101" ELSE
"11101011" WHEN dir_lut ="01110110" ELSE
"11101011" WHEN dir_lut ="01110111" ELSE
"11101100" WHEN dir_lut ="01111000" ELSE
"11101100" WHEN dir_lut ="01111001" ELSE
"11101100" WHEN dir_lut ="01111010" ELSE
"11101100" WHEN dir_lut ="01111011" ELSE
"11101100" WHEN dir_lut ="01111100" ELSE
"11101101" WHEN dir_lut ="01111101" ELSE
"11101101" WHEN dir_lut ="01111110" ELSE
"11101101" WHEN dir_lut ="01111111" ELSE
"11101101" WHEN dir_lut ="10000000" ELSE
"11101101" WHEN dir_lut ="10000001" ELSE
"11101110" WHEN dir_lut ="10000010" ELSE
"11101110" WHEN dir_lut ="10000011" ELSE
"11101110" WHEN dir_lut ="10000100" ELSE
"11101110" WHEN dir_lut ="10000101" ELSE
"11101110" WHEN dir_lut ="10000110" ELSE
"11101111" WHEN dir_lut ="10000111" ELSE
"11101111" WHEN dir_lut ="10001000" ELSE
"11101111" WHEN dir_lut ="10001001" ELSE
"11101111" WHEN dir_lut ="10001010" ELSE
"11101111" WHEN dir_lut ="10001011" ELSE
"11101111" WHEN dir_lut ="10001100" ELSE
"11110000" WHEN dir_lut ="10001101" ELSE
"11110000" WHEN dir_lut ="10001110" ELSE
"11110000" WHEN dir_lut ="10001111" ELSE
"11110000" WHEN dir_lut ="10010000" ELSE
"11110000" WHEN dir_lut ="10010001" ELSE
"11110001" WHEN dir_lut ="10010010" ELSE
"11110001" WHEN dir_lut ="10010011" ELSE
"11110001" WHEN dir_lut ="10010100" ELSE
"11110001" WHEN dir_lut ="10010101" ELSE
"11110001" WHEN dir_lut ="10010110" ELSE
"11110001" WHEN dir_lut ="10010111" ELSE
"11110010" WHEN dir_lut ="10011000" ELSE
"11110010" WHEN dir_lut ="10011001" ELSE
"11110010" WHEN dir_lut ="10011010" ELSE
"11110010" WHEN dir_lut ="10011011" ELSE
"11110010" WHEN dir_lut ="10011100" ELSE
"11110010" WHEN dir_lut ="10011101" ELSE
"11110011" WHEN dir_lut ="10011110" ELSE
"11110011" WHEN dir_lut ="10011111" ELSE
"11110011" WHEN dir_lut ="10100000" ELSE
"11110011" WHEN dir_lut ="10100001" ELSE
"11110011" WHEN dir_lut ="10100010" ELSE
"11110011" WHEN dir_lut ="10100011" ELSE
"11110011" WHEN dir_lut ="10100100" ELSE
"11110100" WHEN dir_lut ="10100101" ELSE
"11110100" WHEN dir_lut ="10100110" ELSE
"11110100" WHEN dir_lut ="10100111" ELSE
"11110100" WHEN dir_lut ="10101000" ELSE
"11110100" WHEN dir_lut ="10101001" ELSE
"11110100" WHEN dir_lut ="10101010" ELSE
"11110101" WHEN dir_lut ="10101011" ELSE
"11110101" WHEN dir_lut ="10101100" ELSE
"11110101" WHEN dir_lut ="10101101" ELSE
"11110101" WHEN dir_lut ="10101110" ELSE
"11110101" WHEN dir_lut ="10101111" ELSE
"11110101" WHEN dir_lut ="10110000" ELSE
"11110101" WHEN dir_lut ="10110001" ELSE
"11110110" WHEN dir_lut ="10110010" ELSE
"11110110" WHEN dir_lut ="10110011" ELSE
"11110110" WHEN dir_lut ="10110100" ELSE
"11110110" WHEN dir_lut ="10110101" ELSE
"11110110" WHEN dir_lut ="10110110" ELSE
"11110110" WHEN dir_lut ="10110111" ELSE
"11110110" WHEN dir_lut ="10111000" ELSE
"11110111" WHEN dir_lut ="10111001" ELSE
"11110111" WHEN dir_lut ="10111010" ELSE
"11110111" WHEN dir_lut ="10111011" ELSE
"11110111" WHEN dir_lut ="10111100" ELSE
"11110111" WHEN dir_lut ="10111101" ELSE
"11110111" WHEN dir_lut ="10111110" ELSE
"11110111" WHEN dir_lut ="10111111" ELSE
"11110111" WHEN dir_lut ="11000000" ELSE
"11111000" WHEN dir_lut ="11000001" ELSE
"11111000" WHEN dir_lut ="11000010" ELSE
"11111000" WHEN dir_lut ="11000011" ELSE
"11111000" WHEN dir_lut ="11000100" ELSE
"11111000" WHEN dir_lut ="11000101" ELSE
"11111000" WHEN dir_lut ="11000110" ELSE
"11111000" WHEN dir_lut ="11000111" ELSE
"11111000" WHEN dir_lut ="11001000" ELSE
"11111001" WHEN dir_lut ="11001001" ELSE
"11111001" WHEN dir_lut ="11001010" ELSE
"11111001" WHEN dir_lut ="11001011" ELSE
"11111001" WHEN dir_lut ="11001100" ELSE
"11111001" WHEN dir_lut ="11001101" ELSE
"11111001" WHEN dir_lut ="11001110" ELSE
"11111001" WHEN dir_lut ="11001111" ELSE
"11111001" WHEN dir_lut ="11010000" ELSE
"11111010" WHEN dir_lut ="11010001" ELSE
"11111010" WHEN dir_lut ="11010010" ELSE
"11111010" WHEN dir_lut ="11010011" ELSE
"11111010" WHEN dir_lut ="11010100" ELSE
"11111010" WHEN dir_lut ="11010101" ELSE
"11111010" WHEN dir_lut ="11010110" ELSE
"11111010" WHEN dir_lut ="11010111" ELSE
"11111010" WHEN dir_lut ="11011000" ELSE
"11111011" WHEN dir_lut ="11011001" ELSE
"11111011" WHEN dir_lut ="11011010" ELSE
"11111011" WHEN dir_lut ="11011011" ELSE
"11111011" WHEN dir_lut ="11011100" ELSE
"11111011" WHEN dir_lut ="11011101" ELSE
"11111011" WHEN dir_lut ="11011110" ELSE
"11111011" WHEN dir_lut ="11011111" ELSE
"11111011" WHEN dir_lut ="11100000" ELSE
"11111011" WHEN dir_lut ="11100001" ELSE
"11111100" WHEN dir_lut ="11100010" ELSE
"11111100" WHEN dir_lut ="11100011" ELSE
"11111100" WHEN dir_lut ="11100100" ELSE
"11111100" WHEN dir_lut ="11100101" ELSE
"11111100" WHEN dir_lut ="11100110" ELSE
"11111100" WHEN dir_lut ="11100111" ELSE
"11111100" WHEN dir_lut ="11101000" ELSE
"11111100" WHEN dir_lut ="11101001" ELSE
"11111100" WHEN dir_lut ="11101010" ELSE
"11111101" WHEN dir_lut ="11101011" ELSE
"11111101" WHEN dir_lut ="11101100" ELSE
"11111101" WHEN dir_lut ="11101101" ELSE
"11111101" WHEN dir_lut ="11101110" ELSE
"11111101" WHEN dir_lut ="11101111" ELSE
"11111101" WHEN dir_lut ="11110000" ELSE
"11111101" WHEN dir_lut ="11110001" ELSE
"11111101" WHEN dir_lut ="11110010" ELSE
"11111101" WHEN dir_lut ="11110011" ELSE
"11111110" WHEN dir_lut ="11110100" ELSE
"11111110" WHEN dir_lut ="11110101" ELSE
"11111110" WHEN dir_lut ="11110110" ELSE
"11111110" WHEN dir_lut ="11110111" ELSE
"11111110" WHEN dir_lut ="11111000" ELSE
"11111110" WHEN dir_lut ="11111001" ELSE
"11111110" WHEN dir_lut ="11111010" ELSE
"11111110" WHEN dir_lut ="11111011" ELSE
"11111110" WHEN dir_lut ="11111100" ELSE
"11111110" WHEN dir_lut ="11111101" ELSE
"11111111" WHEN dir_lut ="11111110" ELSE
"11111111";

end Behavioral;

